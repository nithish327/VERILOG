module moore_overlapping(input clk,rst,in, output reg out);
  reg [2:0]state,next_state;
  parameter s0 = 3'b000,
  s1 = 3'b001,
  s2 = 3'b010,
  s3 = 3'b011,
  s4 = 3'b100;
  always @(posedge clk or posedge rst) begin
    if(rst)
      state <= s0;
    else
      state <= next_state;
  end
    always @(*)begin
      case(state)
        s0:begin
          if (in)
            next_state = s1;
          else
            next_state = s0;
        end
         s1:begin
          if (in)
            next_state = s1;
          else
            next_state = s2;
        end
         s2:begin
          if (in)
            next_state = s3;
          else
            next_state = s0;
        end
         s3:begin
          if (in)
            next_state = s4;
          else
            next_state = s2;
        end
        s4:begin
          if (in)
            next_state = s1;
          else
            next_state = s3;
        end
      endcase
    end
  always @(posedge clk )begin
       if(state==s3 && in)
          out <=1;
        else
          out <=0;
      end
      endmodule
      
