module mod_counter #(parameter n=10)(output reg [3:0]count,
input wire clk, rst
);
always @(posedge clk) begin
    if (rst)
    count <= 4'b0000;
    else if (count == n-1)
    count <= 0;
    else 
    count <= count+1;
end 
endmodule
