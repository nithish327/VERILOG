module tb_full_sub;
  reg a,b,cin;
  wire diff,barrow;
  full_sub dut (.a(a), .b(b), .cin(cin), .diff(diff), .barrow(barrow)); 
  initial begin
    $dumpfile("full_sub.vcd");
    $dumpvars(1,tb_full_sub);
    $monitor("Time =0%t a=%b b=%b cin=%b diff=%b barrow=%b",$time, a, b, cin, diff, barrow);
    a=0; b=0; cin=0;#5
    a=0; b=0; cin=1;#5
    a=0; b=1; cin=0;#5
    a=0; b=1; cin=1;#5
    a=1; b=0; cin=0;#5 
    a=1; b=0; cin=1;#5
    a=1; b=1; cin=0;#5 
    a=1; b=1; cin=1;#5
    $finish;
  end
endmodule
    